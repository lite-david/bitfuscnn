module sim_top ( input wire clk
);

ppu ppu();
  
endmodule