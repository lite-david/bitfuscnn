module sim_top ( input wire clk
);

ppu ppu();
coordinatecomputation coordinatecomputation();
  
endmodule
