module sim_top ( input wire clk
);

ppu ppu();
coordinatecomputation coordinatecomputation();
fusion_unit fusion_unit();
  
endmodule
